
//--------------------------------------------------------------------------------------------------------
// Module  : can_top
// Type    : synthesizable, IP's top
// Standard: Verilog 2001 (IEEE1364-2001)
// Function: CAN bus controller,
//           CAN-TX: buffer input data and send them to CAN bus,
//           CAN-RX: get CAN bus data and output to user
//--------------------------------------------------------------------------------------------------------

module can_top #(
    // local ID parameter
    parameter [10:0] LOCAL_ID      = 11'h456,
    
    // recieve ID filter parameters
    parameter [10:0] RX_ID_SHORT_FILTER = 11'h123,
    parameter [10:0] RX_ID_SHORT_MASK   = 11'h7ff,
    parameter [28:0] RX_ID_LONG_FILTER  = 29'h12345678,
    parameter [28:0] RX_ID_LONG_MASK    = 29'h1fffffff,
    
    // CAN timing parameters
    parameter [15:0] default_c_PTS  = 16'd34,
    parameter [15:0] default_c_PBS1 = 16'd5,
    parameter [15:0] default_c_PBS2 = 16'd10
) (
    input  wire        rstn,      // set to 1 while working
    input  wire        clk,       // system clock
    
    
    // Runtime configuration (optional override for parameters)
    input  wire        cfg_override_en,       // enable runtime configuration
    input  wire [10:0] cfg_local_id,          // runtime TX ID
    input  wire [10:0] cfg_rx_filter_short,   // runtime RX short ID filter
    input  wire [10:0] cfg_rx_mask_short,     // runtime RX short ID mask
    input  wire [28:0] cfg_rx_filter_long,    // runtime RX long ID filter
    input  wire [28:0] cfg_rx_mask_long,      // runtime RX long ID mask
    input  wire [15:0] cfg_c_pts,             // runtime timing: PTS
    input  wire [15:0] cfg_c_pbs1,            // runtime timing: PBS1
    input  wire [15:0] cfg_c_pbs2,            // runtime timing: PBS2
    // CAN TX and RX, connect to external CAN phy (e.g., TJA1050)
    input  wire        can_rx,
    output wire        can_tx,
    
    // user tx-buffer write interface
    input  wire        tx_valid,  // when tx_valid=1 and tx_ready=1, push a data to tx fifo
    output wire        tx_ready,  // whether the tx fifo is available
    input  wire [31:0] tx_data,   // the data to push to tx fifo
    input  wire [ 3:0] tx_len,    // data length (1-4 bytes), if 0 or >4, use 4
    
    // user rx data interface (byte per cycle, unbuffered)
    output reg         rx_valid,  // whether data byte is valid
    output reg         rx_last,   // indicate the last data byte of a packet
    output reg  [ 7:0] rx_data,   // a data byte in the packet
    output reg  [28:0] rx_id,     // the ID of a packet
    output reg         rx_ide     // whether the ID is LONG or SHORT
);



// ---------------------------------------------------------------------------------------------------------------------------------------
//  Runtime configuration selection
// ---------------------------------------------------------------------------------------------------------------------------------------
wire [10:0] local_id_actual        = cfg_override_en ? cfg_local_id        : LOCAL_ID;
wire [10:0] rx_filter_short_actual = cfg_override_en ? cfg_rx_filter_short : RX_ID_SHORT_FILTER;
wire [10:0] rx_mask_short_actual   = cfg_override_en ? cfg_rx_mask_short   : RX_ID_SHORT_MASK;
wire [28:0] rx_filter_long_actual  = cfg_override_en ? cfg_rx_filter_long  : RX_ID_LONG_FILTER;
wire [28:0] rx_mask_long_actual    = cfg_override_en ? cfg_rx_mask_long    : RX_ID_LONG_MASK;
wire [15:0] c_pts_actual           = cfg_override_en ? cfg_c_pts           : default_c_PTS;
wire [15:0] c_pbs1_actual          = cfg_override_en ? cfg_c_pbs1          : default_c_PBS1;
wire [15:0] c_pbs2_actual          = cfg_override_en ? cfg_c_pbs2          : default_c_PBS2;


initial {rx_valid, rx_last, rx_data, rx_id, rx_ide} = 0;

reg         buff_valid = 1'b0;
reg         buff_ready = 1'b0;
wire [31:0] buff_data;
wire [ 3:0] buff_len;   // 缓冲数据长度

reg         pkt_txing = 1'b0;
reg  [31:0] pkt_tx_data = 0;
reg  [ 3:0] pkt_tx_len = 4'd4;  // 发送长度
wire        pkt_tx_done;
wire        pkt_tx_acked;
wire        pkt_rx_valid;
wire [28:0] pkt_rx_id;
wire        pkt_rx_ide;
wire        pkt_rx_rtr;
wire [ 3:0] pkt_rx_len;
wire [63:0] pkt_rx_data;
reg         pkt_rx_ack = 1'b0;

reg         t_rtr_req = 1'b0;
reg         r_rtr_req = 1'b0;
reg  [ 3:0] r_cnt = 4'd0;
reg  [ 3:0] r_len = 4'd0;
reg  [63:0] r_data = 64'h0;
reg  [ 1:0] t_retry_cnt = 2'h0;



// ---------------------------------------------------------------------------------------------------------------------------------------
//  TX buffer
// ---------------------------------------------------------------------------------------------------------------------------------------
localparam DSIZE = 32;
localparam LSIZE = 4;   // 长度字段大小
localparam ASIZE = 2;  //原本是10 我改成2

reg [DSIZE-1:0] buffer [0:((1<<ASIZE)-1)];  // may automatically synthesize to BRAM
reg [LSIZE-1:0] len_buffer [0:((1<<ASIZE)-1)];  // 长度缓冲

reg [ASIZE:0] wptr=0, rptr=0;

wire full  = wptr == {~rptr[ASIZE], rptr[ASIZE-1:0]};
wire empty = wptr == rptr;

assign tx_ready = ~full;

always @ (posedge clk or negedge rstn)
    if(~rstn) begin
        wptr <= 0;
    end else begin
        if(tx_valid & ~full)
            wptr <= wptr + {{ASIZE{1'b0}}, 1'b1};
    end

always @ (posedge clk)
    if(tx_valid & ~full) begin
        buffer[wptr[ASIZE-1:0]] <= tx_data;
        // 存储长度，限制在1-4字节范围
        len_buffer[wptr[ASIZE-1:0]] <= (tx_len == 0 || tx_len > 4) ? 4'd4 : tx_len;
    end

wire            rdready = ~buff_valid | buff_ready;
reg             rdack = 1'b0;
reg [DSIZE-1:0] rddata;
reg [LSIZE-1:0] rdlen;
reg [DSIZE-1:0] keepdata = 0;
reg [LSIZE-1:0] keeplen = 4'd4;
assign buff_data = rdack ? rddata : keepdata;
assign buff_len  = rdack ? rdlen  : keeplen;

always @ (posedge clk or negedge rstn)
    if(~rstn) begin
        buff_valid <= 1'b0;
        rdack <= 1'b0;
        rptr <= 0;
        keepdata <= 0;
        keeplen <= 4'd4;
    end else begin
        buff_valid <= ~empty | ~rdready;
        rdack <= ~empty & rdready;
        if(~empty & rdready)
            rptr <= rptr + {{ASIZE{1'b0}}, 1'b1};
        if(rdack) begin
            keepdata <= rddata;
            keeplen <= rdlen;
        end
    end

always @ (posedge clk) begin
    rddata <= buffer[rptr[ASIZE-1:0]];
    rdlen  <= len_buffer[rptr[ASIZE-1:0]];
end



// ---------------------------------------------------------------------------------------------------------------------------------------
//  CAN packet level controller
// ---------------------------------------------------------------------------------------------------------------------------------------
can_level_packet #(
) u_can_level_packet (
    .rstn            ( rstn             ),
    .clk             ( clk              ),
    
    // Runtime configuration
    .cfg_override_en ( cfg_override_en ),
    .cfg_tx_id       ( local_id_actual ),
    .cfg_c_pts       ( c_pts_actual    ),
    .cfg_c_pbs1      ( c_pbs1_actual   ),
    .cfg_c_pbs2      ( c_pbs2_actual   ),
    
    .can_rx          ( can_rx           ),
    .can_tx          ( can_tx           ),
    
    .tx_start        ( pkt_txing        ),
    .tx_data         ( pkt_tx_data      ),
    .tx_len          ( pkt_tx_len       ),  // 添加长度接口
    .tx_done         ( pkt_tx_done      ),
    .tx_acked        ( pkt_tx_acked     ),
    
    .rx_valid        ( pkt_rx_valid     ),
    .rx_id           ( pkt_rx_id        ),
    .rx_ide          ( pkt_rx_ide       ),
    .rx_rtr          ( pkt_rx_rtr       ),
    .rx_len          ( pkt_rx_len       ),
    .rx_data         ( pkt_rx_data      ),
    .rx_ack          ( pkt_rx_ack       )
);



// ---------------------------------------------------------------------------------------------------------------------------------------
//  RX action
// ---------------------------------------------------------------------------------------------------------------------------------------
always @ (posedge clk or negedge rstn)
    if(~rstn) begin
        pkt_rx_ack <= 1'b0;
        r_rtr_req <= 1'b0;
        r_cnt <= 4'd0;
        r_len <= 4'd0;
        r_data <= 0;
        {rx_valid, rx_last, rx_data, rx_id, rx_ide} <= 0;
    end else begin
        {rx_valid, rx_last, rx_data} <= 0;
        
        pkt_rx_ack <= 1'b0;
        r_rtr_req <= 1'b0;
        
        if(r_cnt>4'd0) begin             // send the data bytes out

            rx_valid <= (r_cnt<=r_len);
            rx_last  <= (r_cnt<=r_len) && (r_cnt==4'd1);
            {rx_data, r_data} <= {r_data, 8'd0};
            r_cnt <= r_cnt - 4'd1;
            
        end else if(pkt_rx_valid) begin  // recieve a new packet
        
            r_len <= pkt_rx_len;             // latches the rx_len
            r_data <= pkt_rx_data;           // latches the rx_data
            
            if(pkt_rx_rtr) begin
                if(~pkt_rx_ide && pkt_rx_id[10:0]==local_id_actual) begin                                           // is a short-ID remote packet, and the ID matches LOCAL_ID
                    pkt_rx_ack <= 1'b1;
                    r_rtr_req <= 1'b1;
                end
            end else if(~pkt_rx_ide) begin                                                                   // is a short-ID data packet
                if( (pkt_rx_id[10:0] & rx_mask_short_actual) == (rx_filter_short_actual & rx_mask_short_actual) ) begin  // ID match
                    pkt_rx_ack <= 1'b1;
                    r_cnt <= 4'd8;
                    rx_id <= pkt_rx_id;
                    rx_ide <= pkt_rx_ide;
                end
            end else begin                                                                                   // is a long-ID data packet
                if( (pkt_rx_id & rx_mask_long_actual) == (rx_filter_long_actual & rx_mask_long_actual) ) begin           // ID match
                    pkt_rx_ack <= 1'b1;
                    r_cnt <= 4'd8;
                    rx_id <= pkt_rx_id;
                    rx_ide <= pkt_rx_ide;
                end
            end
        end
    end



// ---------------------------------------------------------------------------------------------------------------------------------------
//  TX action
// ---------------------------------------------------------------------------------------------------------------------------------------
always @ (posedge clk or negedge rstn)
    if(~rstn) begin
        buff_ready <= 1'b0;
        pkt_tx_data <= 0;
        pkt_tx_len <= 4'd4;
        t_rtr_req <= 1'b0;
        pkt_txing <= 1'b0;
        t_retry_cnt <= 2'd0;
    end else begin
        buff_ready <= 1'b0;

        if(r_rtr_req)
            t_rtr_req <= 1'b1;                   // set t_rtr_req

        if(~pkt_txing) begin
            t_retry_cnt <= 2'd0;
            if(t_rtr_req | buff_valid) begin     // if recieved a remote packet, or tx-buffer data available
                buff_ready <= buff_valid;        // tx-buffer buffer pop, if tx-buffer is available
                t_rtr_req <= 1'b0;               // reset t_rtr_req
                if(buff_valid) begin             // update data from tx-buffer , if tx-buffer is available
                    pkt_tx_data <= buff_data;  // Data should already be left-aligned by caller
                    pkt_tx_len <= buff_len;      // 更新发送长度
                end
                pkt_txing <= 1'b1;
            end
        end else if(pkt_tx_done) begin
            if(pkt_tx_acked || t_retry_cnt==2'd3) begin
                pkt_txing <= 1'b0;
            end else begin
                t_retry_cnt <= t_retry_cnt + 2'd1;
            end
        end
    end


endmodule
